/******************************************************************************
 * (C) Copyright 2021 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * MODULE:      amiq_ofc_defines
 * PROJECT:     Amiq Open-Source Framework for Co-Emulation
 *******************************************************************************/

`ifndef AMIQ_OFC_DEFINES
`define AMIQ_OFC_DEFINES

`define HOSTNAME  "127.0.0.1"
`define PORT      54000
`define END_ITEM  "end_of_test"
`define DELIM     "\n"
`define TIMEOUT   1

`endif
